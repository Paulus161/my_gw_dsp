// designed: Paulus for github

module top ()



endmodule